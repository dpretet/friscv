// copyright damien pretet 2021
// distributed under the mit license
// https://opensource.org/licenses/mit-license.php

`timescale 1 ns / 1 ps
`default_nettype none

module friscv

    #(
    parameter XLEN = 0
    )(
    input         aclk,
    input         aresetn
    );


endmodule

`resetall

