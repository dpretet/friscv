// distributed under the mit license
// https://opensource.org/licenses/mit-license.php

`timescale 1 ns / 1 ps
`default_nettype none

`include "friscv_h.sv"

module friscv_csr

    #(
        parameter RV32E = 0,
        parameter MHART_ID = 0,
        parameter XLEN = 32
    )(
        // clock/reset interface
        input  logic                   aclk,
        input  logic                   aresetn,
        input  logic                   srst,
        // Instruction bus
        input  logic                   valid,
        output logic                   ready,
        input  logic [`INST_BUS_W-1:0] instbus,
        // register source 1 query interface
        output logic [5          -1:0] rs1_addr,
        input  logic [XLEN       -1:0] rs1_val,
        output logic                   rd_wr_en,
        output logic [5          -1:0] rd_wr_addr,
        output logic [XLEN       -1:0] rd_wr_val,
        // External source of CSRs
        input  logic                   ctrl_mepc_wr,
        input  logic [XLEN       -1:0] ctrl_mepc,
        input  logic                   ctrl_mstatus_wr,
        input  logic [XLEN       -1:0] ctrl_mstatus,
        input  logic                   ctrl_mcause_wr,
        input  logic [XLEN       -1:0] ctrl_mcause,
        // status of the processor
        output logic                   ro_trap,
        // CSR shared bus
        output logic [`CSR_SB_W  -1:0] csr_sb
    );

    // ------------------------------------------------------------------------
    // TODO: Ensure CSRRW/CSRRWI read doesn't indude side effect on read if
    //       rd=0 as specified in chapter 9 Zicsr
    // TODO: Print CSR implemented at startup
    // ------------------------------------------------------------------------

    // ------------------------------------------------------------------------
    // Declarations
    // ------------------------------------------------------------------------

    typedef enum logic [1:0] {
        IDLE,
        COMPUTE,
        STORE
    } fsm;

    fsm cfsm;

    // instructions fields
    logic [`OPCODE_W   -1:0] opcode;
    logic [`FUNCT3_W   -1:0] funct3;
    logic [`RS1_W      -1:0] rs1;
    logic [`RD_W       -1:0] rd;
    logic [`ZIMM_W     -1:0] zimm;
    logic [`CSR_W      -1:0] csr;

    logic csr_wren;
    logic csr_rden;
    logic [XLEN-1:0] oldval;
    logic [XLEN-1:0] newval;
    logic [XLEN-1:0] csrs [2**12-1:0];

    logic [`FUNCT3_W -1:0] funct3_r;
    logic [`CSR_W    -1:0] csr_r;
    logic [`ZIMM_W   -1:0] zimm_r;
    logic [5         -1:0] rs1_addr_r;
    logic [XLEN      -1:0] rs1_val_r;

    logic                  ro_write_access;

    // -------------------
    // Machine-level CSRs:
    // -------------------

    // Machine Information Status
    // logic [XLEN-1:0] mvendorid;  // 0xF11    MRO (not implemented)
    // logic [XLEN-1:0] marchid;    // 0xF12    MRO (not implemented)
    // logic [XLEN-1:0] mimpid;     // 0xF13    MRO (not implemented)
    logic [XLEN-1:0] mhartid;       // 0xF14    MRO

    // Machine Trap Status
    logic [XLEN-1:0] mstatus;       // 0x300    MRW
    logic [XLEN-1:0] misa;          // 0x301    MRW
    logic [XLEN-1:0] medeleg;       // 0x302    MRW
    logic [XLEN-1:0] mideleg;       // 0x303    MRW
    logic [XLEN-1:0] mie;           // 0x304    MRW
    logic [XLEN-1:0] mtvec;         // 0x305    MRW
    logic [XLEN-1:0] mcounteren;    // 0x306    MRW

    // Machine Trap Handling
    logic [XLEN-1:0] mscratch;      // 0x340    MRW
    logic [XLEN-1:0] mepc;          // 0x341    MRW
    logic [XLEN-1:0] mcause;        // 0x342    MRW
    logic [XLEN-1:0] mtval;         // 0x343    MRW
    logic [XLEN-1:0] mip;           // 0x344    MRW

    // Machine Memory Protection
    logic [XLEN-1:0] pmpcfg0;       // 0x3A0    MRW
    logic [XLEN-1:0] pmpcfg1;       // 0x3A1    MRW
    logic [XLEN-1:0] pmpcfg2;       // 0x3A2    MRW
    logic [XLEN-1:0] pmpcfg3;       // 0x3A3    MRW
    logic [XLEN-1:0] pmpaddr0;      // 0x3B0    MRW


    // ----------------------
    // Supervisor-level CSRs:
    // ----------------------

    // Supervisor Protection and Translation
    logic [XLEN-1:0] satp;          // 0x180


    // ----------------
    // User-level CSRs:
    // ----------------

    // User Counter/Timers
    logic [XLEN-1:0] cycle;         // 0xC00


    // Logger setup
    svlogger log;
    initial log = new("CSR",
                      `CSR_VERBOSITY,
                      `CSR_ROUTE);

    // ------------------------------------------------------------------------
    // Decompose the instruction bus
    // ------------------------------------------------------------------------

    assign opcode = instbus[`OPCODE +: `OPCODE_W];
    assign funct3 = instbus[`FUNCT3 +: `FUNCT3_W];
    assign rs1    = instbus[`RS1    +: `RS1_W   ];
    assign rd     = instbus[`RD     +: `RD_W    ];
    assign zimm   = instbus[`ZIMM   +: `ZIMM_W  ];
    assign csr    = instbus[`CSR    +: `CSR_W   ];

    assign rs1_addr = rs1;

    // Flags an access which will try to modify a read-only register
    assign ro_write_access = (csr[11:10]==2'b11 && 
                                // only rs1=x0 and these opcodes will be legal
                                ((rs1!=5'b0 &&
                                    (funct3==`CSRRS || funct3==`CSRRC ||
                                    funct3==`CSRRSI || funct3==`CSRRCI)) && 
                                // Any RW opcode is illegal
                                (funct3==`CSRRW && funct3==`CSRRWI))
                             ) ? 1'b1 : 1'b0;

    // ------------------------------------------------------------------------
    // CSR execution machine
    // ------------------------------------------------------------------------

    always @ (posedge aclk or negedge aresetn) begin
        if (aresetn==1'b0) begin
            rd_wr_en <= 1'b0;
            rd_wr_val <= {XLEN{1'b0}};
            ready <= 1'b0;
            csr_wren <= 1'b0;
            newval <= {XLEN{1'b0}};
            funct3_r <= {`FUNCT3_W{1'b0}};
            csr_r <= {`CSR_W{1'b0}};
            zimm_r <= {`ZIMM_W{1'b0}};
            rs1_addr_r <= 5'b0;
            rs1_val_r <= {XLEN{1'b0}};
            rd_wr_addr <= 5'b0;
            ro_trap <= 1'b0;
            cfsm <= IDLE;
        end else if (srst) begin
            rd_wr_en <= 1'b0;
            rd_wr_val <= {XLEN{1'b0}};
            ready <= 1'b0;
            csr_wren <= 1'b0;
            newval <= {XLEN{1'b0}};
            funct3_r <= {`FUNCT3_W{1'b0}};
            csr_r <= {`CSR_W{1'b0}};
            zimm_r <= {`ZIMM_W{1'b0}};
            rs1_addr_r <= 5'b0;
            rs1_val_r <= {XLEN{1'b0}};
            rd_wr_addr <= 5'b0;
            ro_trap <= 1'b0;
            cfsm <= IDLE;
        end else begin

            // Wait for a new instruction
            case(cfsm)

                default: begin

                    csr_wren <= 1'b0;
                    rd_wr_en <= 1'b0;
                    ready <= 1'b1;

                    if (valid) begin
                        if (~ro_write_access) begin
                            ready <= 1'b0;
                            funct3_r <= funct3;
                            csr_r <= csr;
                            zimm_r <= zimm;
                            rs1_addr_r <= rs1;
                            rs1_val_r <= rs1_val;
                            rd_wr_addr <= rd;
                            ro_trap <= 1'b0;
                            cfsm <= COMPUTE;
                        end else begin
                            log.error("Try to write into read-only register");
                            ro_trap <= 1'b1;
                        end
                    end
                end

                // Compute the new CSR value and drive
                // the ISA register
                COMPUTE: begin

                    cfsm <= STORE;

                    // Swap RS1 and CSR
                    if (funct3_r==`CSRRW) begin
                        csr_wren <= 1'b1;
                        rd_wr_en <= 1'b1;
                        rd_wr_val <= oldval;
                        newval <= rs1_val_r;

                    // Save CSR in RS1 and apply a set mask with rs1
                    end else if (funct3_r==`CSRRS) begin
                        rd_wr_en <= 1'b1;
                        rd_wr_val <= oldval;
                        if (rs1_addr_r!=5'b0) begin
                            csr_wren <= 1'b1;
                            newval <= oldval | rs1_val_r;
                        end

                    // Save CSR in RS1 then apply a clear mask fwith rs1
                    end else if (funct3_r==`CSRRC) begin
                        rd_wr_en <= 1'b1;
                        rd_wr_val <= oldval;
                        if (rs1_addr_r!=5'b0) begin
                            csr_wren <= 1'b1;
                            newval <= oldval & rs1_val_r;
                        end

                    // Store CSR in RS1 then set CSR to Zimm
                    end else if (funct3_r==`CSRRWI) begin
                        csr_wren <= 1'b1;
                        rd_wr_en <= 1'b1;
                        rd_wr_val <= oldval;
                        newval <= {{XLEN-5{1'b0}}, zimm_r};

                    // Save CSR in RS1 and apply a set mask with Zimm
                    end else if (funct3_r==`CSRRSI) begin
                        rd_wr_en <= 1'b1;
                        rd_wr_val <= oldval;
                        if (zimm_r!=5'b0) begin
                            csr_wren <= 1'b1;
                            newval <= oldval | {{(XLEN-`ZIMM_W){1'b0}}, zimm_r};
                        end

                    // Save CSR in RS1 and apply a clear mask with Zimm
                    end else if (funct3_r==`CSRRCI) begin
                        rd_wr_en <= 1'b1;
                        rd_wr_val <= oldval;
                        if (zimm_r!=5'b0) begin
                            csr_wren <= 1'b1;
                            newval <= oldval & {{(XLEN-`ZIMM_W){1'b0}}, zimm_r};
                        end

                    end
                end

                // Take time to store new CSR value, handles the
                // RAM behavior according the RAM technology which
                // may be write first / read first. Avoid consecutive
                // CSR instructions to fail
                STORE: begin
                    csr_wren <= 1'b0;
                    rd_wr_en <= 1'b0;
                    if (rd_wr_en==1'b0) begin
                        ready <= 1'b1;
                        cfsm <= IDLE;
                    end
                end
            endcase
        end
    end


    // ------------------------------------------------------------------------
    // CSRs description
    // ------------------------------------------------------------------------

    // HARTID - Read-only
    assign mhartid = MHART_ID;

    // ISA Description: supposed to be RW, is RO in this implementation

    // Supported extensions
    assign misa[0]  = 1'b0;                     // A Atomic extension
    assign misa[1]  = 1'b0;                     // B Tentatively reserved for Bit-Manipulation extension
    assign misa[2]  = 1'b0;                     // C Compressed extension
    assign misa[3]  = 1'b0;                     // D Double-precision floating-point extension
    assign misa[4]  = (RV32E) ? 1'b1 : 1'b0;    // E RV32E base ISA
    assign misa[5]  = 1'b0;                     // F Single-precision floating-point extension
    assign misa[6]  = 1'b0;                     // G Additional standard extensions present
    assign misa[7]  = 1'b0;                     // H Hypervisor extension
    assign misa[8]  = (~RV32E) ? 1'b1 : 1'b0;   // I RV32I/64I/128I base ISA
    assign misa[9]  = 1'b0;                     // J Tentatively reserved for Dynamically Translated Languages extension
    assign misa[10] = 1'b0;                     // K Reserved
    assign misa[11] = 1'b0;                     // L Tentatively reserved for Decimal Floating-Point extension
    assign misa[12] = 1'b0;                     // M Integer Multiply/Divide extension
    assign misa[13] = 1'b0;                     // N User-level interrupts supported
    assign misa[14] = 1'b0;                     // O Reserved
    assign misa[15] = 1'b0;                     // P Tentatively reserved for Packed-SIMD extension
    assign misa[16] = 1'b0;                     // Q Quad-precision floating-point extension
    assign misa[17] = 1'b0;                     // R Reserved
    assign misa[18] = 1'b0;                     // S Supervisor mode implemented
    assign misa[19] = 1'b0;                     // T Tentatively reserved for Transactional Memory extension
    assign misa[20] = 1'b0;                     // U User mode implemented
    assign misa[21] = 1'b0;                     // V Tentatively reserved for Vector extension
    assign misa[22] = 1'b0;                     // W Reserved
    assign misa[23] = 1'b0;                     // X Non-standard extensions present
    assign misa[24] = 1'b0;                     // Y Reserved
    assign misa[25] = 1'b0;                     // Z Reserved


    // MXLEN field encoding
    generate
    if (XLEN==32) begin : MXLEN_32
        assign misa[31:26] = {2'h1, 4'b0};
    end else if (XLEN==64) begin: MXLEN_64
        assign misa[63:26] = {2'h2, 36'b0};
    end else begin: MXLEN_128
        assign misa[127:26] = {2'h3, 100'b0};
    end
    endgenerate

    // TODO: take in account current privilege mode check if rw is applicable

    // MSTATUS (WPRI - Reserved Writes Preserve Values, Reads Ignore Values)
    
    // 31       SD related to XS FS, 0 for the moment
    // 30-23    WPRI
    // 22       TSR Supervisor mode, 0 for the moment
    // 21       TW Timeout Wait, 0 for the moment
    // 20       TVM Virtualization, 0 N/A
    // 19       MXR Virtual Mem, 0 N/A
    // 18       SUM Virtual Mem, 0 N/A
    // 17       MPRV Virtual Mem, 0 N/A
    // 16:15    XS FP, 0 N/A
    // 14:13    FS FP, 0 N/A
    // 12:11    MPP
    // 10:9     WPRI
    // 8        SPP Supervisor mode, 0 for the moment
    // 7        MPIE
    // 6        WPRI
    // 5        SPIE Supervisor mode, 0 for the moment
    // 4        UPIE User mode, 0 for the moment
    // 3        MIE
    // 2        WPRI
    // 1        SIE Supervisor mode, 0 for the moment
    // 0        UIE User mode,  0 for the moment

    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            mstatus <= {XLEN{1'b0}};
        end else if (srst) begin
            mstatus <= {XLEN{1'b0}};
        end else begin
            if (ctrl_mstatus_wr) begin
                mstatus <= {ctrl_mstatus[31], 8'b0, ctrl_mstatus[22:11], 2'b0,
                            ctrl_mstatus[8:7], 1'b0, ctrl_mstatus[5:3], 1'b0,
                            ctrl_mstatus[1:0]};
            end else if (csr_wren) begin
                if (csr_r==12'h300) begin
                    mstatus <= {newval[31], 8'b0, newval[22:11], 2'b0,
                                newval[8:7], 1'b0, newval[5:3], 1'b0,
                                newval[1:0]};
                end
            end
        end
    end 

    // MTVEC (WARL - Write Any Values, Reads Legal Values) 
    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            mtvec <= {XLEN{1'b0}};
        end else if (srst) begin
            mtvec <= {XLEN{1'b0}};
        end else begin
            if (csr_wren) begin
                if (csr_r==12'h305) begin
                    mtvec <= newval;
                end
            end
        end
    end 

    // MSCRATCH
    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            mscratch <= {XLEN{1'b0}};
        end else if (srst) begin
            mscratch <= {XLEN{1'b0}};
        end else begin
            if (csr_wren) begin
                if (csr_r==12'h340) begin
                    mscratch <= newval;
                end
            end
        end
    end 

    // MEPC, only support IALIGN=32
    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            mepc <= {XLEN{1'b0}};
        end else if (srst) begin
            mepc <= {XLEN{1'b0}};
        end else begin
            if (ctrl_mepc_wr) begin
                mepc <= {ctrl_mepc[XLEN-1:2], 2'b0}; 
            end else if (csr_wren) begin
                if (csr_r==12'h341) begin
                    mepc <= {newval[XLEN-1:2], 2'b0};
                end
            end
        end
    end 

    // MCAUSE
    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            mcause <= {XLEN{1'b0}};
        end else if (srst) begin
            mcause <= {XLEN{1'b0}};
        end else begin
            if (ctrl_mcause_wr) begin
                mcause <= ctrl_mcause;
            end else if (csr_wren) begin
                if (csr_r==12'h342) begin
                    mcause <= newval;
                end
            end
        end
    end 

    // MTVAL
    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            mtval <= {XLEN{1'b0}};
        end else if (srst) begin
            mtval <= {XLEN{1'b0}};
        end else begin
            if (csr_wren) begin
                if (csr_r==12'h343) begin
                    mtval <= newval;
                end
            end
        end
    end 


    //////////////////////////////////////////////////////////////////////////
    // Read circuit
    //////////////////////////////////////////////////////////////////////////

    always @ (posedge aclk or negedge aresetn) begin
        if (~aresetn) begin
            oldval <= {XLEN{1'b0}};
        end else if (srst) begin
            oldval <= {XLEN{1'b0}};
        end else begin
            if (cfsm==IDLE && valid) begin
                if (csr==12'h300) begin
                    oldval <= mstatus;
                end else if (csr==12'h301) begin
                    oldval <= misa;
                end else if (csr==12'h305) begin
                    oldval <= mtvec;
                end else if (csr==12'h340) begin
                    oldval <= mscratch;
                end else if (csr==12'h341) begin
                    oldval <= mepc;
                end else if (csr==12'h342) begin
                    oldval <= mcause;
                end else if (csr==12'h343) begin
                    oldval <= mtval;
                end else if (csr==12'hF14) begin
                    oldval <= mhartid;
                end else begin
                    oldval <= {XLEN{1'b0}};
                end
            end
        end
    end


    //////////////////////////////////////////////////////////////////////////
    // CSR Shared bus, for registers used across the processor
    //////////////////////////////////////////////////////////////////////////

    assign csr_sb[`MTVEC+:XLEN] = mtvec;
    assign csr_sb[`MEPC+:XLEN] = mepc;
    assign csr_sb[`MSTATUS+:XLEN] = mstatus;


endmodule

`resetall
