// distributed under the mit license
// https://opensource.org/licenses/mit-license.php

`ifndef FRISCV_DEBUG
`define FRISCV_DEBUG

`define DBG_PC   0
`define DBG_X1   1
`define DBG_X2   2
`define DBG_X3   3
`define DBG_X4   4
`define DBG_X5   5
`define DBG_X6   6
`define DBG_X7   7
`define DBG_X8   8
`define DBG_X9   9
`define DBG_X10  10
`define DBG_X11  11
`define DBG_X12  12
`define DBG_X13  13
`define DBG_X14  14
`define DBG_X15  15
`define DBG_X16  16
`define DBG_X17  17
`define DBG_X18  18
`define DBG_X19  19
`define DBG_X20  20
`define DBG_X21  21
`define DBG_X22  22
`define DBG_X23  23
`define DBG_X24  24
`define DBG_X25  25
`define DBG_X26  26
`define DBG_X27  27
`define DBG_X28  28
`define DBG_X29  29
`define DBG_X30  30
`define DBG_X31  31

`endif
