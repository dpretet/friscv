// distributed under the mit license
// https://opensource.org/licenses/mit-license.php

`ifndef FRISCV_DEBUG
`define FRISCV_DEBUG

`define PC   0
`define X1   1
`define X2   2
`define X3   3
`define X4   4
`define X5   5
`define X6   6
`define X7   7
`define X8   8
`define X9   9
`define X10  10
`define X11  11
`define X12  12
`define X13  13
`define X14  14
`define X15  15
`define X16  16
`define X17  17
`define X18  18
`define X19  19
`define X20  20
`define X21  21
`define X22  22
`define X23  23
`define X24  24
`define X25  25
`define X26  26
`define X27  27
`define X28  28
`define X29  29
`define X30  30
`define X31  31

`endif
