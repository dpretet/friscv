../common/friscv_testbench.sv